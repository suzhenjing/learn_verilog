module su(
    input a
);


endmodule